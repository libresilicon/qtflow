magic
magscale 1 2
timestamp 1522078206793
<< active >>
rect 1600 700 1601 701
rect 1100 600 1101 601
<< contact >>
rect 100 500 300 700
rect 100 900 300 1100
rect 100 1300 300 1500
rect 500 500 700 700
rect 500 900 700 1100
rect 800 1500 801 1501
rect 800 1500 801 1501
rect 700 1500 500 1300
rect 1300 500 1100 700
rect 1300 900 1100 1100
rect 1300 1300 1100 1500
rect 1700 500 1900 700
rect 1800 900 1801 901
rect 200 1200 201 1201
rect 1900 1100 1700 900
rect 1900 1500 1700 1300
rect 2300 700 2500 500
rect 2300 1100 2500 900
rect 2300 1500 2500 1300
rect 2700 1500 2900 1300
rect 2700 1100 2900 900
rect 2700 700 2900 500
rect 1000 100 1200 300
rect 1400 100 1600 300
rect 1800 100 2000 300
<< n_plus_select >>
rect 1400 1600 400 400
rect 2600 1600 3000 400
<< n_well >>
rect 1400 400 0 1600
<< p_plus_select >>
rect 2600 1600 2601 1601
rect 2400 1500 2401 1501
rect 2600 1700 2601 1701
rect 2600 1600 1600 400
rect 0 1600 400 400
<< p_well >>
rect 3000 400 1600 1600
<< poly >>
rect 800 0 2200 400
rect 2100 1700 2101 1701
rect 800 1600 1000 400
rect 2200 400 2000 1600
<< end >>
