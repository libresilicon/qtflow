magic
magscale 1 2
timestamp 1522318414552
<< contact >>
rect 1 8 3 10
rect 1 12 3 14
rect 1 16 3 18
rect 5 8 7 10
rect 5 12 7 14
rect 5 16 7 18
rect 11 8 13 10
rect 11 12 13 14
rect 11 16 13 18
rect 17 8 19 10
rect 17 12 19 14
rect 17 16 19 18
rect 23 8 25 10
rect 23 12 25 14
rect 23 16 25 18
rect 27 8 29 10
rect 27 12 29 14
rect 27 16 29 18
rect 16 2 18 4
rect 12 2 14 4
<< metal1 >>
rect 5 3 5 4
rect 10 5 10 6
rect 18 14 18 15
rect 10 7 20 23
rect 0 0 8 23
rect 30 1 30 1
rect 29 1 29 1
rect 30 21 30 22
rect 22 0 30 23
rect 10 5 20 0
rect 20 0 20 0
<< n_plus_select >>
rect 0 7 4 19
rect 3 4 3 4
rect 26 7 30 19
<< n_well >>
rect 0 7 14 19
<< p_plus_select >>
rect 4 7 14 19
rect 16 7 26 19
<< p_well >>
rect 16 7 30 19
<< poly >>
rect 8 7 10 19
rect 20 7 22 19
rect 8 0 22 7
<< via1 >>
rect 1 20 3 22
rect 5 20 7 22
rect 1 2 3 4
rect 5 2 7 4
rect 23 2 25 4
rect 27 2 29 4
rect 23 20 25 22
rect 27 20 29 22
rect 12 20 14 22
rect 16 20 18 22
<< end >>
