magic
magscale 1 2
timestamp 1521897372782
<< active >>
rect 0 -1400 1400 0
rect 1600 0 3000 -1400
rect 1600 -1000 1601 -999
rect 1100 -1100 1101 -1099
<< contact >>
rect 200 -1200 400 -1000
rect 200 -800 400 -600
rect 200 -400 400 -200
rect 600 -1200 800 -1000
rect 600 -800 800 -600
rect 800 -200 801 -199
rect 800 -200 801 -199
rect 800 -200 600 -400
rect 1200 -1200 1000 -1000
rect 1200 -800 1000 -600
rect 1200 -400 1000 -200
rect 1800 -1200 2000 -1000
rect 1800 -800 1801 -799
rect 200 -500 201 -499
rect 2000 -600 1800 -800
rect 2000 -200 1800 -400
rect 2200 -1000 2400 -1200
rect 2200 -600 2400 -800
rect 2200 -200 2400 -400
rect 2600 -200 2800 -400
rect 2600 -600 2800 -800
rect 2600 -1000 2800 -1200
rect 1000 -1700 1200 -1500
rect 1400 -1700 1600 -1500
rect 1800 -1700 2000 -1500
<< n_well >>
rect 0 0 1400 -1400
<< p_well >>
rect 1600 -1400 3000 0
<< poly >>
rect 800 0 1000 -1400
rect 2000 0 2200 -1400
rect 800 -1800 2200 -1400
<< end >>
